// the register block will be a 32 registers each 32 bits wide

// to address all the blocks in 32 registers, we need to have 4 bits for addressing the register block
module register_block(
    input read_reg_data_1,
    input read_reg_data_2
)

endmodule
